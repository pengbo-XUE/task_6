a   �  a   v   R  o  K  X  �  �      #  7  �  �  �  �  �  �  �  �  �  �     v   FileAndType�   R  �{"baseDir":"C:/Users/Pengb/source/repos/assignment 2 task 6/assignment 2 task 6","file":"obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml","type":"article","sourceDir":"obj/","destinationDir":""}   o  OriginalFileAndType�   K  �{"baseDir":"C:/Users/Pengb/source/repos/assignment 2 task 6/assignment 2 task 6","file":"obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml","type":"article","sourceDir":"obj/","destinationDir":""}   X  KeyJ   �  @~/obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml   �  LocalPathFromRootH     >obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml     LinkToFiles	   #     7  
LinkToUidsI   �  �  �  �  B  ~  �  �    %  E  \  �  �  �  )  H  C   �  9assignment_2_task_6.Models.AddPhoneNumberViewModel.Number;   �  1System.Object.Equals(System.Object,System.Object)D   B  :System.Object.ReferenceEquals(System.Object,System.Object)<   ~  2assignment_2_task_6.Models.AddPhoneNumberViewModel@   �  6System.ComponentModel.DataAnnotations.DisplayAttribute-   �  #System.Object.Equals(System.Object)#     System.Object.GetHashCode   %  System.String    E  System.Object.ToString   \  System.Object$   �  assignment_2_task_6.Models>   �  4System.ComponentModel.DataAnnotations.PhoneAttribute'   �  System.Object.MemberwiseCloneD   )  :assignment_2_task_6.Models.AddPhoneNumberViewModel.Number*   H  System.Object.GetTypeA   �  7System.ComponentModel.DataAnnotations.RequiredAttribute   �  FileLinkSources   �  {}   �  UidLinkSources   �  {}   �  Uids�  �  �[{"name":"assignment_2_task_6.Models.AddPhoneNumberViewModel","file":"obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml"},{"name":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number","file":"obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml"},{"name":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number*","file":"obj/api/assignment_2_task_6.Models.AddPhoneNumberViewModel.yml"}]   �  ManifestProperties   �  {}   �  DocumentType	   �   Zd  .m  {"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.PageViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","items":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"assignment_2_task_6.Models.AddPhoneNumberViewModel","commentId":"T:assignment_2_task_6.Models.AddPhoneNumberViewModel","id":"AddPhoneNumberViewModel","isEii":false,"isExtensionMethod":false,"parent":"assignment_2_task_6.Models","children":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["assignment_2_task_6.Models.AddPhoneNumberViewModel.Number"]},"langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"AddPhoneNumberViewModel","nameWithType":"AddPhoneNumberViewModel","fullName":"assignment_2_task_6.Models.AddPhoneNumberViewModel","type":"Class","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"source/repos/assignment 2 task 6/assignment 2 task 6/Models/ManageViewModels.cs","branch":"master","repo":"https://github.com/pengbo-XUE/Chess_console_v1.git"},"id":"AddPhoneNumberViewModel","path":"Models/ManageViewModels.cs","startLine":60,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["assignment 2 task 6"]},"namespace":"assignment_2_task_6.Models","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"public class AddPhoneNumberViewModel","content.vb":"Public Class AddPhoneNumberViewModel"},"inheritance":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["System.Object"]},"inheritedMembers":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["System.Object.ToString","System.Object.Equals(System.Object)","System.Object.Equals(System.Object,System.Object)","System.Object.ReferenceEquals(System.Object,System.Object)","System.Object.GetHashCode","System.Object.GetType","System.Object.MemberwiseClone"]},"modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","class"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public","Class"]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ItemViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","uid":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number","commentId":"P:assignment_2_task_6.Models.AddPhoneNumberViewModel.Number","id":"Number","isEii":false,"isExtensionMethod":false,"parent":"assignment_2_task_6.Models.AddPhoneNumberViewModel","langs":{"$type":"System.String[], mscorlib","$values":["csharp","vb"]},"name":"Number","nameWithType":"AddPhoneNumberViewModel.Number","fullName":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number","type":"Property","source":{"$type":"Microsoft.DocAsCode.DataContracts.Common.SourceDetail, Microsoft.DocAsCode.DataContracts.Common","remote":{"$type":"Microsoft.DocAsCode.Common.Git.GitDetail, Microsoft.DocAsCode.Common","path":"source/repos/assignment 2 task 6/assignment 2 task 6/Models/ManageViewModels.cs","branch":"master","repo":"https://github.com/pengbo-XUE/Chess_console_v1.git"},"id":"Number","path":"Models/ManageViewModels.cs","startLine":62,"endLine":0,"isExternal":false},"assemblies":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["assignment 2 task 6"]},"namespace":"assignment_2_task_6.Models","syntax":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.SyntaxDetailViewModel, Microsoft.DocAsCode.DataContracts.ManagedReference","content":"[Required]\n[Phone]\n[Display(Name = \"Phone Number\")]\npublic string Number { get; set; }","parameters":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[]},"return":{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.ApiParameter, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.String"},"content.vb":"<Required>\n<Phone>\n<Display(Name:=\"Phone Number\")>\nPublic Property Number As String"},"overload":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number*","attributes":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.AttributeInfo, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.AttributeInfo, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.ComponentModel.DataAnnotations.RequiredAttribute","ctor":"System.ComponentModel.DataAnnotations.RequiredAttribute.#ctor","arguments":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ArgumentInfo, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.AttributeInfo, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.ComponentModel.DataAnnotations.PhoneAttribute","ctor":"System.ComponentModel.DataAnnotations.PhoneAttribute.#ctor","arguments":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ArgumentInfo, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[]}},{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.AttributeInfo, Microsoft.DocAsCode.DataContracts.ManagedReference","type":"System.ComponentModel.DataAnnotations.DisplayAttribute","ctor":"System.ComponentModel.DataAnnotations.DisplayAttribute.#ctor","arguments":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.ArgumentInfo, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[]},"namedArguments":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.ManagedReference.NamedArgumentInfo, Microsoft.DocAsCode.DataContracts.ManagedReference]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.ManagedReference.NamedArgumentInfo, Microsoft.DocAsCode.DataContracts.ManagedReference","name":"Name","type":"System.String","value":"Phone Number"}]}}]},"modifiers.csharp":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["public","get","set"]},"modifiers.vb":{"$type":"System.Collections.Generic.List`1[[System.String, mscorlib]], mscorlib","$values":["Public"]}}]},"references":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"assignment_2_task_6.Models","commentId":"N:assignment_2_task_6.Models","name":"assignment_2_task_6.Models","nameWithType":"assignment_2_task_6.Models","fullName":"assignment_2_task_6.Models"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","commentId":"T:System.Object","parent":"System","isExternal":true,"name":"Object","nameWithType":"Object","fullName":"System.Object"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ToString","commentId":"M:System.Object.ToString","parent":"System.Object","isExternal":true,"name":"ToString()","nameWithType":"Object.ToString()","fullName":"System.Object.ToString()","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ToString","name":"ToString","nameWithType":"Object.ToString","fullName":"System.Object.ToString","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ToString","name":"ToString","nameWithType":"Object.ToString","fullName":"System.Object.ToString","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object)","commentId":"M:System.Object.Equals(System.Object)","parent":"System.Object","isExternal":true,"name":"Equals(Object)","nameWithType":"Object.Equals(Object)","fullName":"System.Object.Equals(System.Object)","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object)","name":"Equals","nameWithType":"Object.Equals","fullName":"System.Object.Equals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object)","name":"Equals","nameWithType":"Object.Equals","fullName":"System.Object.Equals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object,System.Object)","commentId":"M:System.Object.Equals(System.Object,System.Object)","parent":"System.Object","isExternal":true,"name":"Equals(Object, Object)","nameWithType":"Object.Equals(Object, Object)","fullName":"System.Object.Equals(System.Object, System.Object)","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object,System.Object)","name":"Equals","nameWithType":"Object.Equals","fullName":"System.Object.Equals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":", ","nameWithType":", ","fullName":", ","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.Equals(System.Object,System.Object)","name":"Equals","nameWithType":"Object.Equals","fullName":"System.Object.Equals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":", ","nameWithType":", ","fullName":", ","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ReferenceEquals(System.Object,System.Object)","commentId":"M:System.Object.ReferenceEquals(System.Object,System.Object)","parent":"System.Object","isExternal":true,"name":"ReferenceEquals(Object, Object)","nameWithType":"Object.ReferenceEquals(Object, Object)","fullName":"System.Object.ReferenceEquals(System.Object, System.Object)","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ReferenceEquals(System.Object,System.Object)","name":"ReferenceEquals","nameWithType":"Object.ReferenceEquals","fullName":"System.Object.ReferenceEquals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":", ","nameWithType":", ","fullName":", ","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.ReferenceEquals(System.Object,System.Object)","name":"ReferenceEquals","nameWithType":"Object.ReferenceEquals","fullName":"System.Object.ReferenceEquals","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":", ","nameWithType":", ","fullName":", ","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object","name":"Object","nameWithType":"Object","fullName":"System.Object","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetHashCode","commentId":"M:System.Object.GetHashCode","parent":"System.Object","isExternal":true,"name":"GetHashCode()","nameWithType":"Object.GetHashCode()","fullName":"System.Object.GetHashCode()","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetHashCode","name":"GetHashCode","nameWithType":"Object.GetHashCode","fullName":"System.Object.GetHashCode","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetHashCode","name":"GetHashCode","nameWithType":"Object.GetHashCode","fullName":"System.Object.GetHashCode","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetType","commentId":"M:System.Object.GetType","parent":"System.Object","isExternal":true,"name":"GetType()","nameWithType":"Object.GetType()","fullName":"System.Object.GetType()","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetType","name":"GetType","nameWithType":"Object.GetType","fullName":"System.Object.GetType","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.GetType","name":"GetType","nameWithType":"Object.GetType","fullName":"System.Object.GetType","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.MemberwiseClone","commentId":"M:System.Object.MemberwiseClone","parent":"System.Object","isExternal":true,"name":"MemberwiseClone()","nameWithType":"Object.MemberwiseClone()","fullName":"System.Object.MemberwiseClone()","spec.csharp":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.MemberwiseClone","name":"MemberwiseClone","nameWithType":"Object.MemberwiseClone","fullName":"System.Object.MemberwiseClone","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]},"spec.vb":{"$type":"System.Collections.Generic.List`1[[Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common]], mscorlib","$values":[{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.Object.MemberwiseClone","name":"MemberwiseClone","nameWithType":"Object.MemberwiseClone","fullName":"System.Object.MemberwiseClone","isExternal":true},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":"(","nameWithType":"(","fullName":"(","isExternal":false},{"$type":"Microsoft.DocAsCode.DataContracts.Common.SpecViewModel, Microsoft.DocAsCode.DataContracts.Common","name":")","nameWithType":")","fullName":")","isExternal":false}]}},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System","commentId":"N:System","isExternal":true,"name":"System","nameWithType":"System","fullName":"System"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number*","commentId":"Overload:assignment_2_task_6.Models.AddPhoneNumberViewModel.Number","name":"Number","nameWithType":"AddPhoneNumberViewModel.Number","fullName":"assignment_2_task_6.Models.AddPhoneNumberViewModel.Number"},{"$type":"Microsoft.DocAsCode.DataContracts.Common.ReferenceViewModel, Microsoft.DocAsCode.DataContracts.Common","uid":"System.String","commentId":"T:System.String","parent":"System","isExternal":true,"name":"String","nameWithType":"String","fullName":"System.String"}]},"shouldSkipMarkup":false,"_docfxVersion":"2.57.2.0","_systemKeys":{"$type":"System.String[], mscorlib","$values":["uid","isEii","isExtensionMethod","parent","children","href","langs","name","nameWithType","fullName","type","source","documentation","assemblies","namespace","summary","remarks","example","syntax","overridden","overload","exceptions","seealso","see","inheritance","derivedClasses","level","implements","inheritedMembers","extensionMethods","conceptual","platform","attributes","additionalNotes"]}}{   �m  {"$type":"System.Collections.Generic.Dictionary`2[[System.String, mscorlib],[System.Object, mscorlib]], mscorlib"}	   �m   